module Lab4Minterms(
input a,
input b,
input c,
input d,
input e,
input f,
input g,
input h,
input i,
input j,
input k,
output out
);
	assign out = (a&(~b)&(~c)&(~d)&(~e)&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&b&(~c)&(~d)&(~e)&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|(a&b&(~c)&(~d)&(~e)&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|(a&(~b)&c&(~d)&(~e)&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&(~d)&(~e)&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|(a&(~b)&(~c)&d&(~e)&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&b&(~c)&d&(~e)&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&c&d&(~e)&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&(~c)&(~d)&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&b&(~c)&(~d)&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|(a&(~b)&c&(~d)&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&(~d)&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|(a&b&c&(~d)&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&(~c)&d&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|(a&(~b)&(~c)&d&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&b&(~c)&d&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|(a&b&(~c)&d&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&c&d&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|(a&b&c&d&e&(~f)&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&(~c)&(~d)&(~e)&f&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&c&(~d)&(~e)&f&(~g)&(~h)&(~i)&(~j)&(~k))|(a&b&c&(~d)&(~e)&f&(~g)&(~h)&(~i)&(~j)&(~k))|(a&(~b)&(~c)&d&(~e)&f&(~g)&(~h)&(~i)&(~j)&(~k))|(a&b&(~c)&d&(~e)&f&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&d&(~e)&f&(~g)&(~h)&(~i)&(~j)&(~k))|(a&(~b)&(~c)&(~d)&e&f&(~g)&(~h)&(~i)&(~j)&(~k))|(a&(~b)&c&(~d)&e&f&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&(~d)&e&f&(~g)&(~h)&(~i)&(~j)&(~k))|(a&b&c&(~d)&e&f&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&(~c)&d&e&f&(~g)&(~h)&(~i)&(~j)&(~k))|((~a)&b&(~c)&d&e&f&(~g)&(~h)&(~i)&(~j)&(~k))|(a&b&(~c)&d&e&f&(~g)&(~h)&(~i)&(~j)&(~k))|(a&(~b)&(~c)&(~d)&(~e)&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&(~c)&(~d)&(~e)&(~f)&g&(~h)&(~i)&(~j)&(~k))|(a&b&(~c)&(~d)&(~e)&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&(~d)&(~e)&(~f)&g&(~h)&(~i)&(~j)&(~k))|(a&(~b)&(~c)&d&(~e)&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&(~c)&d&(~e)&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&c&d&(~e)&(~f)&g&(~h)&(~i)&(~j)&(~k))|(a&(~b)&c&d&(~e)&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&d&(~e)&(~f)&g&(~h)&(~i)&(~j)&(~k))|(a&b&c&d&(~e)&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&(~c)&(~d)&e&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&(~c)&(~d)&e&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&c&(~d)&e&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&(~d)&e&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&(~c)&d&e&(~f)&g&(~h)&(~i)&(~j)&(~k))|(a&(~b)&(~c)&d&e&(~f)&g&(~h)&(~i)&(~j)&(~k))|(a&b&(~c)&d&e&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&c&d&e&(~f)&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&d&e&(~f)&g&(~h)&(~i)&(~j)&(~k))|(a&b&c&d&e&(~f)&g&(~h)&(~i)&(~j)&(~k))|(a&(~b)&(~c)&(~d)&(~e)&f&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&(~c)&(~d)&(~e)&f&g&(~h)&(~i)&(~j)&(~k))|(a&b&(~c)&(~d)&(~e)&f&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&(~d)&(~e)&f&g&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&(~c)&d&(~e)&f&g&(~h)&(~i)&(~j)&(~k))|(a&(~b)&(~c)&d&(~e)&f&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&(~c)&d&(~e)&f&g&(~h)&(~i)&(~j)&(~k))|((~a)&(~b)&c&d&(~e)&f&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&d&(~e)&f&g&(~h)&(~i)&(~j)&(~k))|(a&(~b)&(~c)&(~d)&e&f&g&(~h)&(~i)&(~j)&(~k))|(a&b&(~c)&(~d)&e&f&g&(~h)&(~i)&(~j)&(~k))|(a&(~b)&c&(~d)&e&f&g&(~h)&(~i)&(~j)&(~k))|((~a)&b&c&(~d)&e&f&g&(~h)&(~i)&(~j)&(~k))|(a&b&c&d&e&f&g&(~h)&(~i)&(~j)&(~k));
endmodule
